CIRCUIT C:\Documents and Settings\All Users\Documents\Softwares\VLSI Softwares\Export Microwind\Example.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
Vclock1 6 0 PULSE(0.00 1.20 20.00N 3.00N 3.00N 20.00N 46.00N)
*
* List of nodes
* "s1" corresponds to n�4
* "clock1" corresponds to n�6
*
* MOS devices
MN1 0 6 4 0 N1  W= 0.36U L= 0.12U
MP1 4 6 1 1 P1  W= 0.36U L= 0.12U
*
C2 1 0  0.764fF
C3 1 0  0.086fF
C4 4 0  0.375fF
C6 6 0  0.176fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.1N 50.00N
* (Pspice)
.PROBE
.END
