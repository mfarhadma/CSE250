* C:\Users\mdfar\OneDrive\Desktop\CSE250\lab\lab 3\Schematic1 lab 3 1.sch

* Schematics Version 9.2
* Tue Jul 27 13:31:58 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic1 lab 3 1.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
